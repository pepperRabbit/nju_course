module my_first_fpga(
	input A,
	input B,
	output F
	);
	
	assign F = ~A&B | A&~B;

endmodule	